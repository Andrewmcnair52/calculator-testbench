`default_nettype none

module test;






initial begin


end








endmodule


